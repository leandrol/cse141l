
module fetch (
	output [2:0] reg_addr1, reg_addr2,
	output [5:0] OPCODE
	);
	
	
endmodule;