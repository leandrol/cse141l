
module ALU (
	input clk,
	input [7:0] IN1, IN2,
	input [5:0] OPCODE,
	output [7:0] result,
	output overflow
	);
	

	
endmodule;