
module fetch (
	input clock,
	input [7:0] program_counter,
	output [8:0] intruction
	);
	
	
	
endmodule;