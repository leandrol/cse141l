
module regfile (
	input clk,
	input [2:0] r_addr1, r_addr2, w_addr,
	input r_or_w,
	output [7:0] data1, data2
	);
	
	
	
endmodule;