module fetch_tb;

	// inputs
	bit clock;
	bit overflow;
	bit bno;
	
	// output
	output [8:0] instruction;
	
endmodule