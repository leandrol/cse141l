
module fetch (
	input clk,
	input [7:0] pc,
	output [2:0] op,
	output [5:0] fields
	);
	
	
endmodule;